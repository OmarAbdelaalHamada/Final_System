module Sys_crtl #(
    parameter FRAME_WIDTH = 8,
    parameter FIFO_DEPTH = 8,
    parameter FIFO_ADDR_WIDTH = $clog2(FIFO_DEPTH),
    parameter ALU_DATA_WIDTH = 16,
    parameter ALU_FUNC_WIDTH = 4,
    parameter REG_FILE_DEPTH = 16,
    parameter REG_FILE_ADDR_WIDTH = $clog2(REG_FILE_DEPTH)
)(
    // Inputs
    input CLK,
    input RST,
    input [ALU_DATA_WIDTH-1:0] ALU_OUT,
    input OUT_VALID,
    input [FRAME_WIDTH-1:0] RdData,
    input RdData_Valid,
    input [FRAME_WIDTH-1:0] RX_P_DATA,
    input RX_P_VLD,
    input FIFO_FULL,

    // Outputs
    output reg [ALU_FUNC_WIDTH-1:0] ALU_FUNC,
    output reg ALU_EN, 
    output reg CLK_EN,
    output reg [REG_FILE_ADDR_WIDTH-1:0] RF_ADDR,
    output reg WrEn,
    output reg RdEn,
    output reg [FRAME_WIDTH-1:0] WrData,
    output reg clk_div_en,
    output reg WR_INC
);

// State Encoding
    
    localparam IDLE           = 4'b0000;
    localparam Rd_Addr        = 4'b0001;
    localparam Rd_Data        = 4'b0011;
    localparam Wr_Addr        = 4'b0010;
    localparam Wr_Data        = 4'b0110;
    localparam Wr_to_RF       = 4'b0111;
    localparam ALU_OP_A       = 4'b0101;
    localparam ALU_OP_B       = 4'b0100;
    localparam ALU_OP_FUNC    = 4'b1100;
    localparam OUT_to_FIFO_1  = 4'b1101;
    localparam OUT_to_FIFO_2  = 4'b1111;
    localparam ALU_NOP_FUNC   = 4'b1110;

// Internal Signals
    reg [3:0] current_state, next_state;
    reg [ALU_DATA_WIDTH-1:0] ALU_OUT_reg;
    reg [REG_FILE_ADDR_WIDTH-1:0] RF_ADDR_reg;
    reg [FRAME_WIDTH-1:0] WrData_reg;

// Internal regs:
// always@(posedge CLK or negedge RST) begin
//     if(!RST) begin
//             ALU_OUT_reg <= 0;
//             RF_ADDR_reg <= 0;
//             WrData_reg <= 0;
//     end
//     else begin

//     end
// end
// State Transition
always @(posedge CLK or negedge RST) begin
    if (!RST) begin
        current_state <= IDLE;
    end else begin
        current_state <= next_state;
    end  
end

// Next State Logic
always @(*) begin
    case (current_state)
        IDLE: begin
           if (RX_P_VLD) begin
                if(RX_P_DATA == 8'hAA) begin 
                    next_state = Wr_Addr;
                end 
                else if(RX_P_DATA == 8'hBB) begin 
                    next_state = Rd_Addr; 
                end
                else if (RX_P_DATA == 8'hCC) begin 
                    next_state = ALU_OP_A; 
                end
                else if (RX_P_DATA == 8'hDD) begin
                    next_state = ALU_NOP_FUNC;
                end
                else begin
                    next_state = IDLE;
                end
            end 
            else begin
                next_state = IDLE;
            end
        end
        Rd_Addr: begin
            if(RX_P_VLD) begin
                next_state = Rd_Data;
            end
            else begin
                next_state = Rd_Addr;
            end
        end
        Rd_Data: begin
            if(RX_P_VLD) begin
                if(RX_P_DATA == 8'hAA) begin 
                    next_state = Wr_Addr;
                end 
                else if(RX_P_DATA == 8'hBB) begin 
                    next_state = Rd_Addr; 
                end
                else if (RX_P_DATA == 8'hCC) begin 
                    next_state = ALU_OP_A; 
                end
                else if (RX_P_DATA == 8'hDD) begin
                    next_state = ALU_NOP_FUNC;
                end
                else begin
                    next_state = IDLE;
                end
            end
            else begin
                next_state = Rd_Data;
            end
        end
        Wr_Addr: begin
            if(RX_P_VLD) begin
                next_state = Wr_Data;
            end
            else begin
                next_state = Wr_Addr;
            end
        end
        Wr_Data: begin
            if(RX_P_VLD) begin
                next_state = Wr_to_RF;
            end
            else begin
                next_state = Wr_Data;
            end
        end
        Wr_to_RF: begin
            if(RX_P_VLD) begin
                if(RX_P_DATA == 8'hAA) begin 
                    next_state = Wr_Addr;
                end 
                else if(RX_P_DATA == 8'hBB) begin 
                    next_state = Rd_Addr; 
                end
                else if (RX_P_DATA == 8'hCC) begin 
                    next_state = ALU_OP_A; 
                end
                else if (RX_P_DATA == 8'hDD) begin
                    next_state = ALU_NOP_FUNC;
                end
                else begin
                    next_state = IDLE;
                end
            end
            else begin
                next_state = Wr_to_RF;
            end
        end
        ALU_OP_A: begin
            if(RX_P_VLD) begin
                next_state = ALU_OP_B;
            end
            else begin
                next_state = ALU_OP_A;
            end
        end
        ALU_OP_B: begin
            if(RX_P_VLD) begin
                next_state = ALU_OP_FUNC;
            end
            else begin
                next_state = ALU_OP_B;
            end
        end
        ALU_OP_FUNC: begin
            if(RX_P_VLD) begin
                next_state = OUT_to_FIFO_1;
            end
            else begin
                next_state = ALU_OP_FUNC;
            end
        end
        OUT_to_FIFO_1: begin
                next_state = OUT_to_FIFO_2;
        end
        OUT_to_FIFO_2: begin
            if(RX_P_VLD) begin
                if(RX_P_DATA == 8'hAA) begin 
                    next_state = Wr_Addr;
                end 
                else if(RX_P_DATA == 8'hBB) begin 
                    next_state = Rd_Addr; 
                end
                else if (RX_P_DATA == 8'hCC) begin 
                    next_state = ALU_OP_A; 
                end
                else if (RX_P_DATA == 8'hDD) begin
                    next_state = ALU_NOP_FUNC;
                end
                else begin
                    next_state = IDLE;
                end
            end
            else begin
                next_state = IDLE;
            end
        end
        ALU_NOP_FUNC: begin
            if(RX_P_VLD) begin
                next_state = OUT_to_FIFO_1;
            end
            else begin
                next_state = ALU_NOP_FUNC;
            end
        end
        default: begin
            next_state = IDLE;
        end
    endcase
end

// Output Logic
always @(*) begin
    ALU_FUNC   = 0;
    ALU_EN     = 0; 
    CLK_EN     = 0;
    RF_ADDR    = 0; 
    WrEn       = 0; 
    RdEn       = 0;
    WrData     = 0; 
    clk_div_en = 1; 
    WR_INC     = 0;
    case (current_state)
        IDLE: begin
            ALU_FUNC   = 0;
            ALU_EN     = 0; 
            CLK_EN     = 0;
            RF_ADDR    = 0; 
            WrEn       = 0; 
            RdEn       = 0;
            WrData     = 0;
            clk_div_en = 1;
        end
        Rd_Addr: begin
            RF_ADDR = RX_P_DATA;
        end
        Rd_Data: begin
            RdEn   = 1;
            clk_div_en = 1;
            if(!FIFO_FULL && RdData_Valid) begin
                WrData = RdData;
                WR_INC = 1;
           end
        end
        Wr_Addr: begin
            RF_ADDR_reg = RX_P_DATA;
            clk_div_en = 1;
        end
        Wr_Data: begin
            WrData_reg = RX_P_DATA;
            clk_div_en = 1;
        end
        Wr_to_RF: begin
            WrEn = 1;
            RF_ADDR = RF_ADDR_reg;
            WrData = WrData_reg;
            clk_div_en = 1;
        end
        ALU_OP_A: begin
            WrEn = 1;
            RF_ADDR = 0;
            WrData = RX_P_DATA;
            clk_div_en = 1;
        end
        ALU_OP_B: begin
            WrEn = 1;
            RF_ADDR = 1;
            WrData = RX_P_DATA;
            clk_div_en = 1;
        end
        ALU_OP_FUNC: begin
            ALU_EN = 1;
            CLK_EN = 1;
            ALU_FUNC = RX_P_DATA[ALU_FUNC_WIDTH-1:0];
            clk_div_en = 1;
        end
        OUT_to_FIFO_1: begin
            ALU_EN = 1;
            CLK_EN = 1;
            clk_div_en = 1;
            ALU_OUT_reg = ALU_OUT;
            if(OUT_VALID && !FIFO_FULL) begin
                WrData  = ALU_OUT_reg[FRAME_WIDTH-1:0];
                WR_INC = 1;
            end
        end
        OUT_to_FIFO_2: begin
            clk_div_en = 1;
            if(!FIFO_FULL) begin
                WrData  = ALU_OUT_reg[2*FRAME_WIDTH-1:FRAME_WIDTH];
                WR_INC = 1;
            end
        end
        ALU_NOP_FUNC: begin
            clk_div_en = 1;
            ALU_EN = 1;
            CLK_EN = 1;
            ALU_FUNC = RX_P_DATA[ALU_FUNC_WIDTH-1:0];
        end
        default: begin
            ALU_FUNC   = 0;
            ALU_EN     = 0; 
            CLK_EN     = 0;
            RF_ADDR    = 0; 
            WrEn       = 0; 
            RdEn       = 0;
            WrData     = 0;
            clk_div_en = 1;
            WR_INC     = 0;
        end
    endcase
end

endmodule